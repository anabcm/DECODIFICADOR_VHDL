LIBRARY ieee;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;    
ENTITY EPROM  is
GENERIC (
BITS: INTEGER:=8;
WORDS: INTEGER:=35
);

PORT ( 
CLKA:IN STD_LOGIC;
addr: IN STD_LOGIC_VECTOR(12 DOWNTO 0);
salida: OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
);
END EPROM;

ARCHITECTURE NARS OF EPROM IS 

TYPE VECTOR_ARRAY IS ARRAY (0 TO WORDS-1) OF STD_LOGIC_VECTOR(13 DOWNTO 0);
CONSTANT memory :vector_array:=(
"00011100000000",--addwf
"00010100000000",--andwf
"00000110000000",--clrf 
"00000100000000",--clrw
"00100100000000",--comf
"00001100000000",--decf
"00101100000000",--decfsz
"00101000000000",---incf
"00111100000000",--infsz
"00010000000000",--iorwf
"00100000000000",--movf
"00000010000000",--movwf
"00000000000000",--nop
"00110100000000",--rlf
"00110000000000",--rrf
"00001000000000",--subwf
"00111000000000",--swapf
"00011000000000",--xorwf
"01000000000000",--bcf
"01010000000000",--bsf
"01100000000000",--btfsc
"01110000000000",--btfss
"11111000000000",--addlw
"11100100000000",--andlw
"10000000000000",--call
"00000001100100",--clrwt
"10100000000000",--goto
"11100000000000",--iorlw
"11000000000000",--movlw
"00000000001001",--retfie
"11010000000000",--retlw
"00000000001000",--return
"00000001100011",--sleep
"11110000000000",--sublw
"11101000000000" --xorlw
);
BEGIN 
PROCESS (addr)
BEGIN 
--IF(CLKA ='1')  THEN
salida<=memory(CONV_INTEGER(addr));
--END IF;
END PROCESS;
end NARS;