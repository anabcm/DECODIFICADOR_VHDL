LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;   
USE IEEE.STD_LOGIC_UNSIGNED.ALL;      
USE IEEE.NUMERIC_BIT.ALL;
ENTITY RAM IS
PORT (
CLKB,RW,CS: in STD_LOGIC;
DIRECCION: in STD_LOGIC_VECTOR(7 DOWN TO 0);
DATAIN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
DATAOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END RAM;
ARCHITECTURE NARQ OF RAM IS
TYPE MEMORIA IS ARRAY (0 TO 511) OF STD_LOGIC(7 DOWNTO O);
SIGNAL RAM:MEMORIA;
BEGIN
PROCESS(CS,RW,CLKB,RAM,DATAIN)
BEGIN
IF(CLKB'EVENT AND CLK='1') THEN
	DATAOUT<=(OTHERS=> 'Z');
	IF (CS='1')THEN
		IF(RW ='0') THEN
			RAM(CONV_INTEGER(DIRECCION))<=DATAIN;
		ELSE
			DATAOUT<=RAM(CONV_INTEGER(DIRECCION));
		END IF;
	END IF;
END IF;
END PROCESS;
END NARQ;