LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECO IS  
PORT (
   CLKA: IN STD_LOGIC;       
   BUS_ENTRA:IN STD_LOGIC_VECTOR(6 DOWNTO 0 );
    SALIDA: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);   
    SD:OUT STD_LOGIC; --DICE SI HAY DIRECCIONAMIENTO INMEDIATO
    ALTA_IMPEDANCIA: OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
);
END DECO;              

ARCHITECTURE NARQ OF DECO IS
BEGIN
PROCESS (CLKA)
VARIABLE CTRL: STD_LOGIC_VECTOR( 1 DOWNTO 0);  --DECODIFICADOR COMPLETO
VARIABLE FROP: STD_LOGIC_VECTOR( 1 DOWNTO 0);   --FILE REGISTER OPERATION
VARIABLE BOFR: STD_LOGIC_VECTOR( 3 DOWNTO 0);   --BYTE ORIENTED FILE REGISTER
VARIABLE LACO: STD_LOGIC_VECTOR( 2 DOWNTO 0);   --BYTE ORIENTED FILE REGISTER  
VARIABLE WR: STD_LOGIC_VECTOR( 1 DOWNTO 0);  --PARA REGISTRO DE TRABAJO         
BEGIN    
CTRL(1):=BUS_ENTRA(6); 
CTRL(0):=BUS_ENTRA(5);   

FROP(1):=BUS_ENTRA(4);
FROP(0):=BUS_ENTRA(3); 
  
BOFR(3):=BUS_ENTRA(4);  
BOFR(2):=BUS_ENTRA(3); 
BOFR(1):=BUS_ENTRA(2);
BOFR(0):=BUS_ENTRA(1); 

LACO(2):=BUS_ENTRA(4); 
LACO(1):=BUS_ENTRA(3); 
LACO(0):=BUS_ENTRA(2); 
     
WR(1):=BUS_ENTRA(4); 
WR(0):=BUS_ENTRA(3); 
IF (CLKA='1') THEN
       ALTA_IMPEDANCIA<="000";--NADIE ESCRIBE EN EL BUS-NI LEE DEL BUS
	CASE CTRL IS
	WHEN "00" =>  SD<='0';
		ALTA_IMPEDANCIA<="001"; --MANEJA UN SALIDA DE F, HABILITA EL MUX MUTANTE Y LE DICE SI PONERSE EN ALTA IMPEDANCIA O NO
		CASE BOFR IS
		    WHEN "0000" =>     --FATA CASO CLRWDT,RETFIE,RETURN,SLEEP
		    		CASE BUS_ENTRA(0) IS
			    		WHEN '0'=>SALIDA<="00001";ALTA_IMPEDANCIA<="111";    --NOP    ALTA IMPEDANCIA NO HACE NADA
			    		WHEN '1'=>SALIDA<="00010";   --MOVWF
		    		END CASE;
		    WHEN "0001" =>
		            CASE BUS_ENTRA(0) IS
			    		WHEN '1'=>SALIDA<="00011";   --CLRF
			    		WHEN '0'=>SALIDA<="00100";ALTA_IMPEDANCIA<="101";   --CLRW   --101 LEE WREG		    		
			    		END CASE;
            WHEN "0010" =>SALIDA<="00101";--SUBWF
            WHEN "0011" =>SALIDA<="00110";--DECF
		    WHEN "0100" =>SALIDA<="00111";--IORWF    
		    WHEN "0101" =>SALIDA<="01000";--ANDWF  
		    WHEN "0110" =>SALIDA<="01001";--XORWF  
		    WHEN "0111" =>SALIDA<="01010";--ADDWF		     
		    WHEN "1000" =>SALIDA<="01011";--MOVF   
		    
		    WHEN "1001" =>SALIDA<="01100";--COMF
		    WHEN "1010" =>SALIDA<="01101";--INCF
		    WHEN "1011" =>SALIDA<="01110";--DECFSZ
            WHEN "1100" =>SALIDA<="01111";--RRF
            WHEN "1101" =>SALIDA<="10000";--RLF  
            
            
            WHEN "1110" =>SALIDA<="10001";--SWAPF
            WHEN "1111" =>SALIDA<="10010";--INCFSZ

		END CASE;
	
	WHEN "01" => SD<='0';ALTA_IMPEDANCIA<="001";--HABILITA EL MUX 	
	      CASE FROP IS
		      WHEN "00"=>SALIDA<="10011";--BCF     
		      WHEN "01"=>SALIDA<="10100";--BSF  
		      WHEN "10"=>SALIDA<="10101";--BTFSC 
		      WHEN "11"=>SALIDA<="10110";--BTFSS   
	      END CASE;	       	
          
	WHEN "10" =>  
		CASE BUS_ENTRA(4) IS
		      WHEN '0'=>SALIDA<="10111";ALTA_IMPEDANCIA<="000";--CALL  --     
		      WHEN '1'=>SALIDA<="11000"; ALTA_IMPEDANCIA<="000";--GOTO         	
		 END CASE;	  
	             SD<='1';

	WHEN "11" =>    SD<='1'; ALTA_IMPEDANCIA<="011";

		CASE WR IS
			WHEN "00"=>SALIDA<="11110"; --MOVLW      si
		END CASE; 
	    CASE LACO IS
	      WHEN "111"=>SALIDA<="11001";--ADDLW si   
	      WHEN "110"=>SALIDA<="11010";--SUBLW  
	      WHEN "101"=>SALIDA<="11011";--XORLW     si
	      WHEN "100"=> 
		      CASE BUS_ENTRA(1) is
			      WHEN '0'=>SALIDA<="11100";--IORLW  
			      WHEN '1'=>SALIDA<="11101";--ANDLW
		      END CASE;	 
	      END CASE;
	          
	WHEN OTHERS => SALIDA<="00000";  
    END CASE;
END IF;
END PROCESS;
END NARQ;

