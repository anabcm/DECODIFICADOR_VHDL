--MUXMUTANTE                 
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADDMUX IS  
PORT (      
RESET,CLKB,CLKD: IN STD_LOGIC;
DIRADD:IN STD_LOGIC_VECTOR(6 DOWNTO 0); 		 --DIRECTO
INDADD:IN STD_LOGIC_VECTOR(7 DOWNTO 0);           --INDIRECTO     
BUSD:INOUT STD_LOGIC_VECTOR(7 DOWNTO 0); 
STATIN:IN STD_LOGIC_VECTOR(2 DOWNTO 0);           --ENTRADA A STATUS
DIRECCION: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);      --DIRECCION GENERADA
E: IN STD_LOGIC;            
E_RAM:OUT STD_LOGIC;
ALTA_IMPEDANCIA: IN STD_LOGIC_VECTOR(2 DOWNTO 0)
);
END ADDMUX;


ARCHITECTURE NARQ OF ADDMUX IS    
BEGIN  
   
PROCESS (CLKB,CLKD,STATIN)     --CALCULA LA DIRECCION  a buscar en RAM     
VARIABLE STATUS: STD_LOGIC_VECTOR(7 DOWNTO 0);         --!irp!rp1!rp0!  to!pd!z!dc!c
VARIABLE FSR: STD_LOGIC_VECTOR(7 DOWNTO 0);        
VARIABLE PCL: STD_LOGIC_VECTOR(7 DOWNTO 0);  
BEGIN     
--IF(   STATIN 'EVENT ) THEN  
 --      STATUS(2 DOWNTO 0)<=STATUSIN;
--END IF;
IF(ALTA_IMPEDANCIA="001") THEN

	IF(CLKB 'EVENT AND CLKB='1') THEN  
		BUSD<="ZZZZZZZZ"; 
		E_RAM<='0';

		CASE DIRADD IS
		WHEN "0000000" => --DIRECCINAMIENTO INDIRECTO 
		           DIRECCION(7 DOWNTO 0)<=INDADD(7 DOWNTO 0);
		           DIRECCION(8)<=STATUS(7);   
		WHEN "0000010" =>DIRECCION<="000000010";--PCL      
		WHEN "0000011"=>DIRECCION<="000000011";--STATUS
		WHEN "0000100"=>DIRECCION<="000000100";--FSR
		WHEN OTHERS =>    
		           DIRECCION(6 DOWNTO 0)<=DIRADD(6 DOWNTO 0);
		           DIRECCION(7)<=STATUS(5);   
		           DIRECCION(7)<=STATUS(6);
		             E_RAM<='1';
		END CASE;   
	END IF;
	
	IF(STATIN 'EVENT AND STATIN='1') THEN                      
	           STATUS(2):=STATIN (2);      
	           STATUS(1):=STATIN (1);     
	           STATUS(0):=STATIN (0);  
	 END IF;                            
	 IF(CLKD 'EVENT AND CLKD='1') THEN 
	 	E_RAM<='0';
	    CASE DIRADD IS
	    WHEN "0000010" =>PCL:=BUSD;--PCL      
		WHEN "0000011"=>STATUS:=BUSD;--STATUS
		WHEN "0000100"=>FSR:=BUSD;--FSR 
		WHEN OTHERS => E_RAM<='1';
        END CASE;
	 
	 END IF;
ELSE
	  	BUSD<="ZZZZZZZZ";
END IF;

END PROCESS; 


END NARQ;                                                                     
