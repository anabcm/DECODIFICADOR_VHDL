--INTRUCTION REG
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY INS_REG IS  
PORT (     
PROGRAM_BUS:IN STD_LOGIC_VECTOR(13 DOWNTO 0);
DIRECT_ADDR:OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
DECO_BUS: OUT STD_LOGIC_VECTOR(6 DOWNTO 0); 
BIT_OPERA: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
CONS:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END INS_REG;

ARCHITECTURE NARQ OF INS_REG IS
BEGIN
PROCESS (PROGRAM_BUS)     
	BEGIN  
	DIRECT_ADDR<=PROGRAM_BUS(6 DOWNTO 0);
	DECO_BUS<=PROGRAM_BUS(13 DOWNTO 7);
	BIT_OPERA<=PROGRAM_BUS(11 DOWNTO 9);
	CONS<=PROGRAM_BUS(7 DOWNTO 0);		
	END PROCESS;
END NARQ;

