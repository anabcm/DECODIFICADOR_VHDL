LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY  WREG IS
PORT( 
ENTRA: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
SALE: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);   
ALTA_IMPEDANCIA: IN STD_LOGIC_VECTOR(2 DOWNTO 0);

CLKD: IN STD_LOGIC
);
END WREG;

ARCHITECTURE NARQ OF WREG IS
BEGIN     

PROCESS (CLKD,ALTA_IMPEDANCIA)
	BEGIN    
	IF ALTA_IMPEDANCIA="011"  THEN
	IF CLKD='1'  AND CLKD'EVENT   THEN
	SALE<=ENTRA;
	END IF;  
	ELSE    ENTRA<="ZZZZZZZZ";
	END IF;

END PROCESS;
END NARQ;           